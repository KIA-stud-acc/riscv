module top();
 riscv_ps rvps();
 instrMem im();
 dataMem  dm();
endmodule